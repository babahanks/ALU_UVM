//`include "alu_top.sv"
//`include "alu.sv"
`include "alu_top.sv"